class out_data;
	logic [9:0] b10_data; 
	logic start_out;
endclass : out_data
