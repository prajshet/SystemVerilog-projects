// 32 bit Table for CRC generation
function [31:0] crcTable;
    input [7:0] data;
    begin
    case(data)
		0: crcTable=32'h00000000;
        1: crcTable=32'h77073096;
        2: crcTable=32'hEE0E612C;
        3: crcTable=32'h990951BA;
        4: crcTable=32'h076DC419;
        5: crcTable=32'h706AF48F;
        6: crcTable=32'hE963A535;
        7: crcTable=32'h9E6495A3;
        8: crcTable=32'h0EDB8832;
        9: crcTable=32'h79DCB8A4;
        10: crcTable=32'hE0D5E91E;
        11: crcTable=32'h97D2D988;
        12: crcTable=32'h09B64C2B;
        13: crcTable=32'h7EB17CBD;
        14: crcTable=32'hE7B82D07;
        15: crcTable=32'h90BF1D91;
        16: crcTable=32'h1DB71064;
        17: crcTable=32'h6AB020F2;
        18: crcTable=32'hF3B97148;
        19: crcTable=32'h84BE41DE;
        20: crcTable=32'h1ADAD47D;
        21: crcTable=32'h6DDDE4EB;
        22: crcTable=32'hF4D4B551;
        23: crcTable=32'h83D385C7;
        24: crcTable=32'h136C9856;
        25: crcTable=32'h646BA8C0;
        26: crcTable=32'hFD62F97A;
        27: crcTable=32'h8A65C9EC;
        28: crcTable=32'h14015C4F;
        29: crcTable=32'h63066CD9;
        30: crcTable=32'hFA0F3D63;
        31: crcTable=32'h8D080DF5;
        32: crcTable=32'h3B6E20C8;
        33: crcTable=32'h4C69105E;
        34: crcTable=32'hD56041E4;
        35: crcTable=32'hA2677172;
        36: crcTable=32'h3C03E4D1;
        37: crcTable=32'h4B04D447;
        38: crcTable=32'hD20D85FD;
        39: crcTable=32'hA50AB56B;
        40: crcTable=32'h35B5A8FA;
        41: crcTable=32'h42B2986C;
        42: crcTable=32'hDBBBC9D6;
        43: crcTable=32'hACBCF940;
        44: crcTable=32'h32D86CE3;
        45: crcTable=32'h45DF5C75;
        46: crcTable=32'hDCD60DCF;
        47: crcTable=32'hABD13D59;
        48: crcTable=32'h26D930AC;
        49: crcTable=32'h51DE003A;
        50: crcTable=32'hC8D75180;
        51: crcTable=32'hBFD06116;
        52: crcTable=32'h21B4F4B5;
        53: crcTable=32'h56B3C423;
        54: crcTable=32'hCFBA9599;
        55: crcTable=32'hB8BDA50F;
        56: crcTable=32'h2802B89E;
        57: crcTable=32'h5F058808;
        58: crcTable=32'hC60CD9B2;
        59: crcTable=32'hB10BE924;
        60: crcTable=32'h2F6F7C87;
        61: crcTable=32'h58684C11;
        62: crcTable=32'hC1611DAB;
        63: crcTable=32'hB6662D3D;
        64: crcTable=32'h76DC4190;
        65: crcTable=32'h01DB7106;
        66: crcTable=32'h98D220BC;
        67: crcTable=32'hEFD5102A;
        68: crcTable=32'h71B18589;
        69: crcTable=32'h06B6B51F;
        70: crcTable=32'h9FBFE4A5;
        71: crcTable=32'hE8B8D433;
        72: crcTable=32'h7807C9A2;
        73: crcTable=32'h0F00F934;
        74: crcTable=32'h9609A88E;
        75: crcTable=32'hE10E9818;
        76: crcTable=32'h7F6A0DBB;
        77: crcTable=32'h086D3D2D;
        78: crcTable=32'h91646C97;
        79: crcTable=32'hE6635C01;
        80: crcTable=32'h6B6B51F4;
        81: crcTable=32'h1C6C6162;
        82: crcTable=32'h856530D8;
        83: crcTable=32'hF262004E;
        84: crcTable=32'h6C0695ED;
        85: crcTable=32'h1B01A57B;
        86: crcTable=32'h8208F4C1;
        87: crcTable=32'hF50FC457;
        88: crcTable=32'h65B0D9C6;
        89: crcTable=32'h12B7E950;
        90: crcTable=32'h8BBEB8EA;
        91: crcTable=32'hFCB9887C;
        92: crcTable=32'h62DD1DDF;
        93: crcTable=32'h15DA2D49;
        94: crcTable=32'h8CD37CF3;
        95: crcTable=32'hFBD44C65;
        96: crcTable=32'h4DB26158;
        97: crcTable=32'h3AB551CE;
        98: crcTable=32'hA3BC0074;
        99: crcTable=32'hD4BB30E2;
        100: crcTable=32'h4ADFA541;
        101: crcTable=32'h3DD895D7;
        102: crcTable=32'hA4D1C46D;
        103: crcTable=32'hD3D6F4FB;
        104: crcTable=32'h4369E96A;
        105: crcTable=32'h346ED9FC;
        106: crcTable=32'hAD678846;
        107: crcTable=32'hDA60B8D0;
        108: crcTable=32'h44042D73;
        109: crcTable=32'h33031DE5;
        110: crcTable=32'hAA0A4C5F;
        111: crcTable=32'hDD0D7CC9;
        112: crcTable=32'h5005713C;
        113: crcTable=32'h270241AA;
        114: crcTable=32'hBE0B1010;
        115: crcTable=32'hC90C2086;
        116: crcTable=32'h5768B525;
        117: crcTable=32'h206F85B3;
        118: crcTable=32'hB966D409;
        119: crcTable=32'hCE61E49F;
        120: crcTable=32'h5EDEF90E;
        121: crcTable=32'h29D9C998;
        122: crcTable=32'hB0D09822;
        123: crcTable=32'hC7D7A8B4;
        124: crcTable=32'h59B33D17;
        125: crcTable=32'h2EB40D81;
        126: crcTable=32'hB7BD5C3B;
        127: crcTable=32'hC0BA6CAD;
        128: crcTable=32'hEDB88320;
        129: crcTable=32'h9ABFB3B6;
        130: crcTable=32'h03B6E20C;
        131: crcTable=32'h74B1D29A;
        132: crcTable=32'hEAD54739;
        133: crcTable=32'h9DD277AF;
        134: crcTable=32'h04DB2615;
        135: crcTable=32'h73DC1683;
        136: crcTable=32'hE3630B12;
        137: crcTable=32'h94643B84;
        138: crcTable=32'h0D6D6A3E;
        139: crcTable=32'h7A6A5AA8;
        140: crcTable=32'hE40ECF0B;
        141: crcTable=32'h9309FF9D;
        142: crcTable=32'h0A00AE27;
        143: crcTable=32'h7D079EB1;
        144: crcTable=32'hF00F9344;
        145: crcTable=32'h8708A3D2;
        146: crcTable=32'h1E01F268;
        147: crcTable=32'h6906C2FE;
        148: crcTable=32'hF762575D;
        149: crcTable=32'h806567CB;
        150: crcTable=32'h196C3671;
        151: crcTable=32'h6E6B06E7;
        152: crcTable=32'hFED41B76;
        153: crcTable=32'h89D32BE0;
        154: crcTable=32'h10DA7A5A;
        155: crcTable=32'h67DD4ACC;
        156: crcTable=32'hF9B9DF6F;
        157: crcTable=32'h8EBEEFF9;
        158: crcTable=32'h17B7BE43;
        159: crcTable=32'h60B08ED5;
        160: crcTable=32'hD6D6A3E8;
        161: crcTable=32'hA1D1937E;
        162: crcTable=32'h38D8C2C4;
        163: crcTable=32'h4FDFF252;
        164: crcTable=32'hD1BB67F1;
        165: crcTable=32'hA6BC5767;
        166: crcTable=32'h3FB506DD;
        167: crcTable=32'h48B2364B;
        168: crcTable=32'hD80D2BDA;
        169: crcTable=32'hAF0A1B4C;
        170: crcTable=32'h36034AF6;
        171: crcTable=32'h41047A60;
        172: crcTable=32'hDF60EFC3;
        173: crcTable=32'hA867DF55;
        174: crcTable=32'h316E8EEF;
        175: crcTable=32'h4669BE79;
        176: crcTable=32'hCB61B38C;
        177: crcTable=32'hBC66831A;
        178: crcTable=32'h256FD2A0;
        179: crcTable=32'h5268E236;
        180: crcTable=32'hCC0C7795;
        181: crcTable=32'hBB0B4703;
        182: crcTable=32'h220216B9;
        183: crcTable=32'h5505262F;
        184: crcTable=32'hC5BA3BBE;
        185: crcTable=32'hB2BD0B28;
        186: crcTable=32'h2BB45A92;
        187: crcTable=32'h5CB36A04;
        188: crcTable=32'hC2D7FFA7;
        189: crcTable=32'hB5D0CF31;
        190: crcTable=32'h2CD99E8B;
        191: crcTable=32'h5BDEAE1D;
        192: crcTable=32'h9B64C2B0;
        193: crcTable=32'hEC63F226;
        194: crcTable=32'h756AA39C;
        195: crcTable=32'h026D930A;
        196: crcTable=32'h9C0906A9;
        197: crcTable=32'hEB0E363F;
        198: crcTable=32'h72076785;
        199: crcTable=32'h05005713;
        200: crcTable=32'h95BF4A82;
        201: crcTable=32'hE2B87A14;
        202: crcTable=32'h7BB12BAE;
        203: crcTable=32'h0CB61B38;
        204: crcTable=32'h92D28E9B;
        205: crcTable=32'hE5D5BE0D;
        206: crcTable=32'h7CDCEFB7;
        207: crcTable=32'h0BDBDF21;
        208: crcTable=32'h86D3D2D4;
        209: crcTable=32'hF1D4E242;
        210: crcTable=32'h68DDB3F8;
        211: crcTable=32'h1FDA836E;
        212: crcTable=32'h81BE16CD;
        213: crcTable=32'hF6B9265B;
        214: crcTable=32'h6FB077E1;
        215: crcTable=32'h18B74777;
        216: crcTable=32'h88085AE6;
        217: crcTable=32'hFF0F6A70;
        218: crcTable=32'h66063BCA;
        219: crcTable=32'h11010B5C;
        220: crcTable=32'h8F659EFF;
        221: crcTable=32'hF862AE69;
        222: crcTable=32'h616BFFD3;
        223: crcTable=32'h166CCF45;
        224: crcTable=32'hA00AE278;
        225: crcTable=32'hD70DD2EE;
        226: crcTable=32'h4E048354;
        227: crcTable=32'h3903B3C2;
        228: crcTable=32'hA7672661;
        229: crcTable=32'hD06016F7;
        230: crcTable=32'h4969474D;
        231: crcTable=32'h3E6E77DB;
        232: crcTable=32'hAED16A4A;
        233: crcTable=32'hD9D65ADC;
        234: crcTable=32'h40DF0B66;
        235: crcTable=32'h37D83BF0;
        236: crcTable=32'hA9BCAE53;
        237: crcTable=32'hDEBB9EC5;
        238: crcTable=32'h47B2CF7F;
        239: crcTable=32'h30B5FFE9;
        240: crcTable=32'hBDBDF21C;
        241: crcTable=32'hCABAC28A;
        242: crcTable=32'h53B39330;
        243: crcTable=32'h24B4A3A6;
        244: crcTable=32'hBAD03605;
        245: crcTable=32'hCDD70693;
        246: crcTable=32'h54DE5729;
        247: crcTable=32'h23D967BF;
        248: crcTable=32'hB3667A2E;
        249: crcTable=32'hC4614AB8;
        250: crcTable=32'h5D681B02;
        251: crcTable=32'h2A6F2B94;
        252: crcTable=32'hB40BBE37;
        253: crcTable=32'hC30C8EA1;
        254: crcTable=32'h5A05DF1B;
        255: crcTable=32'h2D02EF8D;
	endcase
    end
endfunction