// message object from ref_b5 encoder model
class en_data;
logic [9:0] enco;
logic  enco_start;
endclass:en_data
