// message object from input monitor 

class in_data ;

logic [8:0] si_data; //din
logic start_dis ;  // start in
//logic end_dis;
endclass : in_data
